/*
my_hdmi_device

Copyright (C) 2021  Hirosh Dabui <hirosh@dabui.de>

Permission to use, copy, modify, and/or distribute this software for any
purpose with or without fee is hereby granted, provided that the above
copyright notice and this permission notice appear in all copies.

THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
*/
module chip_balls (
    input clk_25mhz,
    output [3:0] gpdi_dp,
    output [7:0] led
);

  reg [7:0] vga_red;
  reg [7:0] vga_blue;
  reg [7:0] vga_green;

  reg vga_hsync;
  reg vga_vsync;
  reg vga_blank;

  localparam SYSTEM_CLK_MHZ = 25;
  localparam DDR_HDMI_TRANSFER = 1;

  // calculate video timings
  localparam x_res = 1280;
  localparam y_res = 720;
  /* localparam x_res             = 640; */
  /* localparam y_res             = 480; */
  localparam frame_rate = 60;

  `include "video_timings.v"

  // clock generator
  wire clk_locked;
  wire [3:0] clocks;

  ecp5pll #(
      .in_hz  (SYSTEM_CLK_MHZ * 1e6),
      .out0_hz(pixel_f * (DDR_HDMI_TRANSFER ? 5 : 10)),
      .out1_hz(pixel_f)
  ) ecp5pll_inst (
      .clk_i (clk_25mhz),
      .clk_o (clocks),
      .locked(clk_locked)
  );

  wire tmds_clk = clocks[0];
  wire pclk = clocks[1];

  wire [10:0] hcnt;
  wire [10:0] vcnt;
  wire hcycle;
  wire vcycle;
  wire hsync;
  wire vsync;
  wire blank;

  my_vga_clk_generator  /*
    //  one of my monitor dislikes autogenerated calculated values
    // just use default vga values in my_vga_clk_generator.vh
    #(
      .VPOL( 1 ),
      .HPOL( 1 ),
      .FRAME_RATE( frame_rate ),
      .VBP( vsync_back_porch ),
      .VFP( vsync_front_porch ),
      .VSLEN( vsync_pulse_width ),
      .VACTIVE( y_res ),
      .HBP( hsync_back_porch ),
      .HFP( hsync_front_porch ),
      .HSLEN( hsync_pulse_width ),
      .HACTIVE( x_res )
    )
    */
  my_vga_clk_generator_i (
      .pclk(pclk),
      .out_hcnt(hcnt),
      .out_vcnt(vcnt),
      .out_hsync(hsync),
      .out_vsync(vsync),
      .out_blank(blank),
      .reset_n(1'b1)
  );

  reg [31:0] frame_cnt = 0;
  wire new_frame = (vcnt == 0 && hcnt == 0);
  wire fps = frame_cnt == 59;
  reg toogle;
  always @(posedge pclk) begin
    if (new_frame) frame_cnt <= fps ? 0 : frame_cnt + 1;
    //toogle <= fps ? !toogle : toogle;
    toogle <= toogle ^ fps;
  end

  assign led = {8{toogle}};

  localparam N = 35;
  wire [N-1:0] draw_ball;
  //reg [N-1:0] in_opposite = 0;
  genvar i;
  generate
    for (i = 0; i < N; i = i + 1) begin : gen_ball
      ball #(
          .START_X(i * 10 % x_res),
          .START_Y(i * 10 % y_res),
          .DELTA_X(1 + (i) % 4),
          .DELTA_Y(1 + (i) % 4),
          .BALL_WIDTH(10 + i % 100),
          .BALL_HEIGHT(10 + i % 100),
          .X_RES(x_res),
          .Y_RES(y_res)
      ) ball_i (
          .clk(pclk),
          .i_vcnt(vcnt),
          .i_hcnt(hcnt),
          //.in_opposite(in_opposite[i]),
          .i_opposite(1'b0),
          .o_draw(draw_ball[i])
      );
    end
  endgenerate
  /////////////////////
  wire [15:0] lfsr;
  wire draw_stars = hcnt >= 0 && hcnt < 256 && vcnt >= 0 && vcnt < 256;
  wire star_object = (&lfsr[15:6] & draw_stars);
  LFSR #(16'b1_0000_0000_1011, 0) lfsr_i (
      pclk,
      1'b0,
      draw_stars,
      lfsr
  );

  wire [15:0] lfsr1;
  wire draw_stars1 = hcnt >= 256 && hcnt < 512 && vcnt >= 0 && vcnt < 256;
  wire star_object1 = (&lfsr1[15:6] & draw_stars1);
  LFSR #(16'b1000000001011, 0) lfsr_i1 (
      pclk,
      1'b0,
      draw_stars1,
      lfsr1
  );

  wire [15:0] lfsr2;
  wire draw_stars2 = hcnt >= 512 && hcnt < (512 + 256) && vcnt >= 0 && vcnt < 256;
  wire star_object2 = (&lfsr2[15:6] & draw_stars2);
  LFSR #(16'b1000000001011, 0) lfsr_i2 (
      pclk,
      1'b0,
      draw_stars2,
      lfsr2
  );

  //////

  wire [15:0] lfsr3;
  wire draw_stars3 = hcnt >= 0 && hcnt < 256 && vcnt >= 224 && vcnt < 480;
  wire star_object3 = (&lfsr3[15:6] & draw_stars3);
  LFSR #(16'b1000000001011, 0) lfsr_i3 (
      pclk,
      1'b0,
      draw_stars3,
      lfsr3
  );

  wire [15:0] lfsr4;
  wire draw_stars4 = hcnt >= 256 && hcnt < 512 && vcnt >= 224 && vcnt < 480;
  wire star_object4 = (&lfsr4[15:6] & draw_stars4);
  LFSR #(16'b1000000001011, 0) lfsr_i4 (
      pclk,
      1'b0,
      draw_stars4,
      lfsr4
  );

  wire [15:0] lfsr5;
  wire draw_stars5 = hcnt >= 512 && hcnt < (512 + 256) && vcnt >= 224 && vcnt < 480;
  wire star_object5 = (&lfsr5[15:6] & draw_stars5);
  LFSR #(16'b1000000001011, 0) lfsr_i5 (
      pclk,
      1'b0,
      draw_stars5,
      lfsr5
  );

  wire stars = star_object  | star_object1 |
     star_object2 | star_object3 |
     star_object4 | star_object5;
  /////////////////////
  wire [7:0] W = {8{hcnt[7:0] == vcnt[7:0]}};
  wire [7:0] A = {8{hcnt[7:5] == 3'h2 && vcnt[7:5] == 3'h2}};
  wire [7:0] vga_red_test = ({hcnt[5:0] & {6{vcnt[4:3] == ~hcnt[4:3]}}, 2'b00} | W) & ~A;
  wire [7:0] vga_green_test = (hcnt[7:0] & {8{vcnt[6]}} | W) & ~A;
  wire [7:0] vga_blue_test = vcnt[7:0] | W | A;

  always @(posedge pclk) begin
    vga_blank <= blank;
    vga_hsync <= hsync;
    vga_vsync <= vsync;

    if (~blank) begin
      vga_red   <= vga_red_test>>1   | (stars | |draw_ball[10:0] | |draw_ball[20:11] | (&vcnt[4:0]|&hcnt[4:0]) ? 8'hff : 8'h0);
      vga_green <= vga_green_test >> 1 | (stars | |draw_ball[20:11] ? 8'hff : 8'h0);
      vga_blue  <= vga_blue_test>>1  | (stars | |draw_ball[34:21] | (&vcnt[4:0]|&hcnt[4:0]) ? 8'hff : 8'h0);
    end else begin
      vga_red   <= 8'h0;
      vga_blue  <= 8'h0;
      vga_green <= 8'h0;
    end
  end

  localparam OUT_TMDS_MSB = DDR_HDMI_TRANSFER ? 1 : 0;
  wire [OUT_TMDS_MSB:0] out_tmds_red;
  wire [OUT_TMDS_MSB:0] out_tmds_green;
  wire [OUT_TMDS_MSB:0] out_tmds_blue;
  wire [OUT_TMDS_MSB:0] out_tmds_clk;

  hdmi_device #(
      .DDR_ENABLED(DDR_HDMI_TRANSFER)
  ) hdmi_device_i (
      pclk,
      tmds_clk,

      vga_red,
      vga_green,
      vga_blue,

      vga_blank,
      vga_vsync,
      vga_hsync,

      out_tmds_red,
      out_tmds_green,
      out_tmds_blue,
      out_tmds_clk
  );

  /* ulx3s can SDR and DDR */
  generate
    if (DDR_HDMI_TRANSFER) begin
      ODDRX1F ddr0_clock (
          .D0(out_tmds_clk   [0] ),
          .D1(out_tmds_clk   [1] ),
          .Q(gpdi_dp[3]),
          .SCLK(tmds_clk),
          .RST(0)
      );
      ODDRX1F ddr0_red (
          .D0(out_tmds_red   [0] ),
          .D1(out_tmds_red   [1] ),
          .Q(gpdi_dp[2]),
          .SCLK(tmds_clk),
          .RST(0)
      );
      ODDRX1F ddr0_green (
          .D0(out_tmds_green[0]),
          .D1(out_tmds_green[1]),
          .Q(gpdi_dp[1]),
          .SCLK(tmds_clk),
          .RST(0)
      );
      ODDRX1F ddr0_blue (
          .D0(out_tmds_blue[0]),
          .D1(out_tmds_blue[1]),
          .Q(gpdi_dp[0]),
          .SCLK(tmds_clk),
          .RST(0)
      );
    end else begin
      assign gpdi_dp[3] = out_tmds_clk;
      assign gpdi_dp[2] = out_tmds_red;
      assign gpdi_dp[1] = out_tmds_green;
      assign gpdi_dp[0] = out_tmds_blue;
    end
  endgenerate

endmodule
